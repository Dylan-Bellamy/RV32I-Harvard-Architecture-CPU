-- megafunction wizard: %RAM: 1-port%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altsyncram 

-- ============================================================
-- File Name: system_memory.vhd
-- Megafunction Name(s):
-- 			altsyncram
--
-- Simulation library Files(s):
-- 			altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THis FILE!
--
-- 13.0.1 Build 232 06/12/2013 SP 1 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2013 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


library ieee;
use ieee.std_logic_1164.all;

library altera_mf;
use altera_mf.all;

entity system_memory is
	port
	(
		address		: in std_logic_vector (5 downto 0);
		clock		: in std_logic  := '1';
		data		: in std_logic_vector (31 downto 0);
		wren		: in std_logic ;
		q		: out std_logic_vector (31 downto 0)
	);
end system_memory;


architecture SYN of system_memory is

	signal sub_wire0	: std_logic_vector (31 downto 0);



	component altsyncram
	generic (
		clock_enable_input_a		: string;
		clock_enable_output_a		: string;
		init_file		: string;
		intended_device_family		: string;
		lpm_hint		: string;
		lpm_type		: string;
		numwords_a		: natural;
		operation_mode		: string;
		outdata_aclr_a		: string;
		outdata_reg_a		: string;
		power_up_uninitialized		: string;
		widthad_a		: natural;
		width_a		: natural;
		width_byteena_a		: natural
	);
	port (
			address_a	: in std_logic_vector (5 downto 0);
			clock0	: in std_logic ;
			data_a	: in std_logic_vector (31 downto 0);
			wren_a	: in std_logic ;
			q_a	: out std_logic_vector (31 downto 0)
	);
	end component;

begin
	q    <= sub_wire0(31 downto 0);

	altsyncram_component : altsyncram
	generic MAP (
		clock_enable_input_a => "BYPASS",
		clock_enable_output_a => "BYPASS",
		init_file => "system_memory.mif",
		intended_device_family => "Cyclone II",
		lpm_hint => "ENABLE_RUNTIME_MOD=NO",
		lpm_type => "altsyncram",
		numwords_a => 64,
		operation_mode => "SINGLE_port",
		outdata_aclr_a => "NONE",
		outdata_reg_a => "CLOCK0",
		power_up_uninitialized => "FALSE",
		widthad_a => 6,
		width_a => 32,
		width_byteena_a => 1
	)
	port MAP (
		address_a => address,
		clock0 => clock,
		data_a => data,
		wren_a => wren,
		q_a => sub_wire0
	);



end SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: ADDRESSSTALL_A NUMERIC "0"
-- Retrieval info: PRIVATE: AclrAddr NUMERIC "0"
-- Retrieval info: PRIVATE: AclrByte NUMERIC "0"
-- Retrieval info: PRIVATE: AclrData NUMERIC "0"
-- Retrieval info: PRIVATE: Aclroutput NUMERIC "0"
-- Retrieval info: PRIVATE: BYTE_ENABLE NUMERIC "0"
-- Retrieval info: PRIVATE: BYTE_SIZE NUMERIC "8"
-- Retrieval info: PRIVATE: BlankMemory NUMERIC "0"
-- Retrieval info: PRIVATE: CLOCK_ENABLE_inPUT_A NUMERIC "0"
-- Retrieval info: PRIVATE: CLOCK_ENABLE_outPUT_A NUMERIC "0"
-- Retrieval info: PRIVATE: Clken NUMERIC "0"
-- Retrieval info: PRIVATE: DataBusSeparated NUMERIC "1"
-- Retrieval info: PRIVATE: IMPLEMENT_in_LES NUMERIC "0"
-- Retrieval info: PRIVATE: inIT_FILE_LAYout string "port_A"
-- Retrieval info: PRIVATE: inIT_TO_SIM_X NUMERIC "0"
-- Retrieval info: PRIVATE: inTendED_DEVICE_FAMILY string "Cyclone II"
-- Retrieval info: PRIVATE: JTAG_ENABLED NUMERIC "0"
-- Retrieval info: PRIVATE: JTAG_ID string "NONE"
-- Retrieval info: PRIVATE: MAXIMUM_DEPTH NUMERIC "0"
-- Retrieval info: PRIVATE: MIFfilename string "system_memory.mif"
-- Retrieval info: PRIVATE: NUMWORDS_A NUMERIC "64"
-- Retrieval info: PRIVATE: RAM_BLOCK_TYPE NUMERIC "0"
-- Retrieval info: PRIVATE: READ_DURinG_WRITE_MODE_port_A NUMERIC "3"
-- Retrieval info: PRIVATE: RegAddr NUMERIC "1"
-- Retrieval info: PRIVATE: RegData NUMERIC "1"
-- Retrieval info: PRIVATE: Regoutput NUMERIC "1"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX string "0"
-- Retrieval info: PRIVATE: SingleClock NUMERIC "1"
-- Retrieval info: PRIVATE: useDQRAM NUMERIC "1"
-- Retrieval info: PRIVATE: WRCONTROL_ACLR_A NUMERIC "0"
-- Retrieval info: PRIVATE: WidthAddr NUMERIC "6"
-- Retrieval info: PRIVATE: WidthData NUMERIC "32"
-- Retrieval info: PRIVATE: rden NUMERIC "0"
-- Retrieval info: library: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: CLOCK_ENABLE_inPUT_A string "BYPASS"
-- Retrieval info: CONSTANT: CLOCK_ENABLE_outPUT_A string "BYPASS"
-- Retrieval info: CONSTANT: inIT_FILE string "system_memory.mif"
-- Retrieval info: CONSTANT: inTendED_DEVICE_FAMILY string "Cyclone II"
-- Retrieval info: CONSTANT: LPM_HinT string "ENABLE_RUNTIME_MOD=NO"
-- Retrieval info: CONSTANT: LPM_TYPE string "altsyncram"
-- Retrieval info: CONSTANT: NUMWORDS_A NUMERIC "64"
-- Retrieval info: CONSTANT: OPERATION_MODE string "SinGLE_port"
-- Retrieval info: CONSTANT: outDATA_ACLR_A string "NONE"
-- Retrieval info: CONSTANT: outDATA_REG_A string "CLOCK0"
-- Retrieval info: CONSTANT: POWER_UP_UNinITIALIZED string "FALSE"
-- Retrieval info: CONSTANT: WIDTHAD_A NUMERIC "6"
-- Retrieval info: CONSTANT: WIDTH_A NUMERIC "32"
-- Retrieval info: CONSTANT: WIDTH_BYTEENA_A NUMERIC "1"
-- Retrieval info: useD_port: address 0 0 6 0 inPUT NODEFVAL "address[5..0]"
-- Retrieval info: useD_port: clock 0 0 0 0 inPUT VCC "clock"
-- Retrieval info: useD_port: data 0 0 32 0 inPUT NODEFVAL "data[31..0]"
-- Retrieval info: useD_port: q 0 0 32 0 outPUT NODEFVAL "q[31..0]"
-- Retrieval info: useD_port: wren 0 0 0 0 inPUT NODEFVAL "wren"
-- Retrieval info: CONNECT: @address_a 0 0 6 0 address 0 0 6 0
-- Retrieval info: CONNECT: @clock0 0 0 0 0 clock 0 0 0 0
-- Retrieval info: CONNECT: @data_a 0 0 32 0 data 0 0 32 0
-- Retrieval info: CONNECT: @wren_a 0 0 0 0 wren 0 0 0 0
-- Retrieval info: CONNECT: q 0 0 32 0 @q_a 0 0 32 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL system_memory.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL system_memory.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL system_memory.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL system_memory.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL system_memory_inst.vhd FALSE
-- Retrieval info: LIB_FILE: altera_mf
